module test #(
    p = 10
) (
    input  a,
    output b
);
endmodule