module dcs_packet_rx_v2 #(
    parameter pDataWidth = 20,
    parameter pBaud = 115_200
    )(
    input iClk
    );
endmodule