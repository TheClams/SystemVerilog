module arithm_op_port #(
	pq_symbols = 4
	)(
	output logic [pq_symbols*4-1:0] name
	);
endmodule