package my_pkg;

   localparam int WIDTH = 16;
   localparam int WIDTH_P1 = WIDTH+1;
   //
   localparam logic [1:0] VECT2B = 2'b10;

endpackage
