module simple();endmodule