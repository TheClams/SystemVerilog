module m();
    logic a;
endmodule