function void f();
    int x=0;
    `uvm_fatal("x","y")
    x++;
endfunction