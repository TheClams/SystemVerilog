module m1 (



input  wire signed a10, aa10,
output wire signed b10, bb10,
inout wire signed c10, cc10,

input  wire unsigned a11, aa11,
output wire unsigned b11, bb11,
inout wire unsigned c11, cc11,

output reg dump
);

endmodule