module m1 (
input a, 
input reg [1:0] b,
input signed c,
input wire d
);
endmodule
