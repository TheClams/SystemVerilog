module m3();
    generate
    endgenerate
endmodule