module a();
logic aaaa [bw];
logic aaaaaa[bw];
logic aaaaa[bw];
logic aaa[bw];
endmodule