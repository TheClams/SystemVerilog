module dcs_packet_rx_v2 #(
pDataWidth = 20,
pBaud = 115_200
)(
input iClk
);
endmodule