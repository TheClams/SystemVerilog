that one is fake "certainly//"? // but me
first comment
/*comment*/
second
//comment
///comment
/*//*/
big comment
/*comment
comment*/
that one is fake "certainly//"?
may and that one "nope" //comment
multi fake "/*not me*/"
int/**/x=5;