module a();
    logic aaaa  [bw]   ;
    logic aaaaaa[bw]   ;
    logic aa           ;
    logic aaaaa [bw][4];
    logic aaa   [bw]   ;
endmodule