class myclass extends baseclass;

    extern function func1 ();
    extern virtual function func2 ();

endclass

